/**
* This file would contain all the definitions needed for the test bench
* 	--RedNdu
*/

/** ALU Operations timing */ 

// BIT ENCODING: 001X XXXD DDDD SSSS Siii iiii iiii iiii
`define CYCLES_ADDI 1
`define CYCLES_SUBI 1
`define CYCLES_ANDI 1
`define CYCLES_ORI  1
`define CYCLES_XORI 1
`define CYCLES_SHLI 1
`define CYCLES_SHRI 1

// BIT ENCODING: 0011 011D DDDD SSSS STTT TTZZ ZZZZ ZXXX
`define CYCLES_ADD  1
`define CYCLES_SUB  1
`define CYCLES_MULT 1
`define CYCLES_AND  1
`define CYCLES_OR   1
`define CYCLES_XOR  1
`define CYCLES_SHR  1
`define CYCLES_SHL  1

// BIT ENCODING: 0011 101D DDDD SSSS STTT TTZZ ZZZZ ZZXX
`define CYCLES_FADD  1
`define CYCLES_FSUB  1
`define CYCLES_FMULT 1
`define CYCLES_FDIV  1

// BIT ENCODING: 0001 00XD DDDD ZZii iiii iiii iiii iiii
`define CYCLES_LIH  1
`define CYCLES_LIL  1

// BIT ENCODING: 0XXX XXXD DDDD SSSS STTT TTZZ ZZZZ EEEE 
`define CYCLES_VADD  1
`define CYCLES_VSUB  1
`define CYCLES_VMULT 1
`define CYCLES_VDIV	 1
`define CYCLES_VDOT  1
`define CYCLES_VDOTA 1

// BIT ENCODING: 0100 101D DDDD TTTT TZZZ ZZZi iZZZ ZZZZ
`define CYCLES_VINDX  1

// BIT ENCODING: 0100 11XD DDDD TTTT TZZZ ZZZZ ZZZZ EEEE
`define CYCLES_VREDUCE 1
`define CYCLES_VSPLAT  1

// BIT ENCODING: 0101 000D DDDD SSSS S112 2334 4ZZZ EEEE
`define CYCLES_VSWIZZLE  1

// BIT ENCODING: 0101 000D DDDD SSSS S112 2334 4ZZZ EEEE
`define CYCLES_VSADD  1
`define CYCLES_VSMULT 1
`define CYCLES_VSSUB  1
`define CYCLES_VSDIV  1

// BIT ENCODING: 0101 101D DDDD SSSS STTT TTCC CCCZ EEEE
`define CYCLES_VSMA 1

